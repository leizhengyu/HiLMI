module LMI#(parameter WR_NUM=4,RD_NUM=4)(
input 


);

